* On-die Decoupling circuit for Z90B (VDDQ to VSSQ)
* Includes VDDQ-VSSQ decoupling for an individual signal such as DQ0-15, LDQS_t/c, UDQS_t/c, UDM or LDM.
* This subcircuit should be added across the IBIS DQ, DM or DQS model's [Pullup Reference] and [Pulldown Reference]
* nodes as in the following Spice example:

******************************************************************************************************
*x_decouple vddq_die vcc_die vssq_die gnd z90b_ondie_decoupling_perdq

*b_dq1 vccq_die vssq_die PAD_DQ1 IN_DQ1 ENOUT RCVR_OUT_DQ1 vccq_die vssq_die
*+ file='z90b.ibs' model='DQ_34_2666' typ=typ power=off buffer=3 interpol=1 ramp_fwf=2 ramp_rwf=2
*+ rm_tail_rwf=default rm_tail_fwf=default
*+ rm_dly_rwf=default rm_dly_fwf=default
******************************************************************************************************


.subckt z90b_ondie_decoupling_perdq vddq_die vcc_die vssq_die ref
x1 vddq_die ref vcc_die ref vssq_die ref z90b_cfat_perdq


**********************************************************
** STATE-SPACE REALIZATION               
** IN SPICE LANGUAGE
** This file is automatically generated  
**********************************************************
** Created: 06-Apr-2017 by IdEM R2012 (8.0.6)
**********************************************************


**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt z90b_cfat_perdq
+  a_1 b_1 
+  a_2 b_2 
+  a_3 b_3 
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+001
GC_1_1 b_1 NI_1 NS_1 0 6.2330481876482144e-002
GC_1_2 b_1 NI_1 NS_2 0 1.4713375097713654e-003
GC_1_3 b_1 NI_1 NS_3 0 5.3402244987502156e-005
GC_1_4 b_1 NI_1 NS_4 0 2.9916990101003390e-004
GC_1_5 b_1 NI_1 NS_5 0 6.3605358032491108e-009
GC_1_6 b_1 NI_1 NS_6 0 8.2886093490834400e-006
GC_1_7 b_1 NI_1 NS_7 0 -4.6276292791965212e-013
GC_1_8 b_1 NI_1 NS_8 0 -6.3862148638194715e-012
GC_1_9 b_1 NI_1 NS_9 0 6.1064222637401668e-002
GC_1_10 b_1 NI_1 NS_10 0 5.1474876326707171e-004
GC_1_11 b_1 NI_1 NS_11 0 -5.5536131048513680e-005
GC_1_12 b_1 NI_1 NS_12 0 -5.9272904883043206e-004
GC_1_13 b_1 NI_1 NS_13 0 -5.3323109299307199e-009
GC_1_14 b_1 NI_1 NS_14 0 5.6127000392586824e-008
GC_1_15 b_1 NI_1 NS_15 0 -9.5370055414972298e-013
GC_1_16 b_1 NI_1 NS_16 0 -7.4859516679077225e-012
GC_1_17 b_1 NI_1 NS_17 0 6.0384528734901126e-002
GC_1_18 b_1 NI_1 NS_18 0 1.4214648197082016e-003
GC_1_19 b_1 NI_1 NS_19 0 4.0023396818858168e-005
GC_1_20 b_1 NI_1 NS_20 0 2.9788583204761539e-004
GC_1_21 b_1 NI_1 NS_21 0 1.8301436759807446e-009
GC_1_22 b_1 NI_1 NS_22 0 -8.3444029837943225e-006
GC_1_23 b_1 NI_1 NS_23 0 1.7536923220494038e-012
GC_1_24 b_1 NI_1 NS_24 0 1.3827429167130989e-011
GD_1_1 b_1 NI_1 NA_1 0 -2.2213701341043574e-001
GD_1_2 b_1 NI_1 NA_2 0 6.0303899466092374e-002
GD_1_3 b_1 NI_1 NA_3 0 5.9921072993829420e-002
*
* Port 2
VI_2 a_2 NI_2 0
RI_2 NI_2 b_2 5.0000000000000000e+001
GC_2_1 b_2 NI_2 NS_1 0 6.1089596134556882e-002
GC_2_2 b_2 NI_2 NS_2 0 5.1273388778624450e-004
GC_2_3 b_2 NI_2 NS_3 0 -5.5557793331426699e-005
GC_2_4 b_2 NI_2 NS_4 0 -5.9272919069189084e-004
GC_2_5 b_2 NI_2 NS_5 0 -5.2417620455036903e-009
GC_2_6 b_2 NI_2 NS_6 0 5.7141036703498026e-008
GC_2_7 b_2 NI_2 NS_7 0 3.2378255712926917e-014
GC_2_8 b_2 NI_2 NS_8 0 9.8152539411647279e-014
GC_2_9 b_2 NI_2 NS_9 0 6.4630999006333512e-002
GC_2_10 b_2 NI_2 NS_10 0 1.6048392606398305e-003
GC_2_11 b_2 NI_2 NS_11 0 1.1890366224678413e-004
GC_2_12 b_2 NI_2 NS_12 0 1.1741287261270675e-003
GC_2_13 b_2 NI_2 NS_13 0 6.5794287495325816e-009
GC_2_14 b_2 NI_2 NS_14 0 1.6035145301151459e-009
GC_2_15 b_2 NI_2 NS_15 0 2.7588828263331523e-012
GC_2_16 b_2 NI_2 NS_16 0 -1.5113333502281194e-012
GC_2_17 b_2 NI_2 NS_17 0 6.2261420630156425e-002
GC_2_18 b_2 NI_2 NS_18 0 4.0917509344954434e-004
GC_2_19 b_2 NI_2 NS_19 0 -5.1215362769534793e-005
GC_2_20 b_2 NI_2 NS_20 0 -5.9020141819952335e-004
GC_2_21 b_2 NI_2 NS_21 0 9.8939063062027746e-010
GC_2_22 b_2 NI_2 NS_22 0 -5.8864369645544587e-008
GC_2_23 b_2 NI_2 NS_23 0 -2.4581234500619735e-012
GC_2_24 b_2 NI_2 NS_24 0 1.3692150323449172e-012
GD_2_1 b_2 NI_2 NA_1 0 6.0267759327233689e-002
GD_2_2 b_2 NI_2 NA_2 0 -2.2111458036981552e-001
GD_2_3 b_2 NI_2 NA_3 0 6.1129898132990003e-002
*
* Port 3
VI_3 a_3 NI_3 0
RI_3 NI_3 b_3 5.0000000000000000e+001
GC_3_1 b_3 NI_3 NS_1 0 6.0409961489978112e-002
GC_3_2 b_3 NI_3 NS_2 0 1.4195048779714994e-003
GC_3_3 b_3 NI_3 NS_3 0 4.0010708122684294e-005
GC_3_4 b_3 NI_3 NS_4 0 2.9788574955973461e-004
GC_3_5 b_3 NI_3 NS_5 0 1.7483522291849174e-009
GC_3_6 b_3 NI_3 NS_6 0 -8.3454142388175917e-006
GC_3_7 b_3 NI_3 NS_7 0 7.6758629823654600e-013
GC_3_8 b_3 NI_3 NS_8 0 6.2438973845733984e-012
GC_3_9 b_3 NI_3 NS_9 0 6.2261423594070088e-002
GC_3_10 b_3 NI_3 NS_10 0 4.0918718196107889e-004
GC_3_11 b_3 NI_3 NS_11 0 -5.1220058734527679e-005
GC_3_12 b_3 NI_3 NS_12 0 -5.9020143266096895e-004
GC_3_13 b_3 NI_3 NS_13 0 1.0749945975704755e-009
GC_3_14 b_3 NI_3 NS_14 0 -5.7850253149727278e-008
GC_3_15 b_3 NI_3 NS_15 0 -1.4720530023322780e-012
GC_3_16 b_3 NI_3 NS_16 0 8.9533199293688142e-012
GC_3_17 b_3 NI_3 NS_17 0 6.1282913495898844e-002
GC_3_18 b_3 NI_3 NS_18 0 1.3752541256966866e-003
GC_3_19 b_3 NI_3 NS_19 0 4.1774874932237504e-005
GC_3_20 b_3 NI_3 NS_20 0 2.9664008114032447e-004
GC_3_21 b_3 NI_3 NS_21 0 -9.8275348283841851e-010
GC_3_22 b_3 NI_3 NS_22 0 8.4026980527323762e-006
GC_3_23 b_3 NI_3 NS_23 0 1.0371174134860775e-012
GC_3_24 b_3 NI_3 NS_24 0 -1.5240513888925418e-011
GD_3_1 b_3 NI_3 NA_1 0 5.9884368428755691e-002
GD_3_2 b_3 NI_3 NA_2 0 6.1129862128178378e-002
GD_3_3 b_3 NI_3 NA_3 0 -2.2173952402741595e-001
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+000
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-002
*
* Impinging wave, port 2
RA_2 NA_2 0 3.5355339059327378e+000
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 b_2 2.0000000000000000e-002
*
* Impinging wave, port 3
RA_3 NA_3 0 3.5355339059327378e+000
FA_3 0 NA_3 VI_3 1.0
GA_3 0 NA_3 a_3 b_3 2.0000000000000000e-002
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-013
RS_1 NS_1 0 2.9502412466187273e+000
GS_1_1 0 NS_1 NA_1 0 6.6452709208363170e-001
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-013
RS_2 NS_2 0 9.7963963778649585e+000
GS_2_1 0 NS_2 NA_1 0 6.6452709208363170e-001
*
* Real pole n. 3
CS_3 NS_3 0 9.9999999999999998e-013
RS_3 NS_3 0 3.6187013423789601e+001
GS_3_1 0 NS_3 NA_1 0 6.6452709208363170e-001
*
* Real pole n. 4
CS_4 NS_4 0 9.9999999999999998e-013
RS_4 NS_4 0 4.6620502512561899e+002
GS_4_1 0 NS_4 NA_1 0 6.6452709208363170e-001
*
* Real pole n. 5
CS_5 NS_5 0 9.9999999999999998e-013
RS_5 NS_5 0 3.0454843143654548e+003
GS_5_1 0 NS_5 NA_1 0 6.6452709208363170e-001
*
* Real pole n. 6
CS_6 NS_6 0 9.9999999999999998e-013
RS_6 NS_6 0 4.2483511278785496e+004
GS_6_1 0 NS_6 NA_1 0 6.6452709208363170e-001
*
* Real pole n. 7
CS_7 NS_7 0 9.9999999999999998e-013
RS_7 NS_7 0 1.7479012563424539e+007
GS_7_1 0 NS_7 NA_1 0 6.6452709208363170e-001
*
* Real pole n. 8
CS_8 NS_8 0 9.9999999999999998e-013
RS_8 NS_8 0 7.6442948626474559e+007
GS_8_1 0 NS_8 NA_1 0 6.6452709208363170e-001
*
* Real pole n. 9
CS_9 NS_9 0 9.9999999999999998e-013
RS_9 NS_9 0 2.9502412466187273e+000
GS_9_2 0 NS_9 NA_2 0 6.6452709208363170e-001
*
* Real pole n. 10
CS_10 NS_10 0 9.9999999999999998e-013
RS_10 NS_10 0 9.7963963778649585e+000
GS_10_2 0 NS_10 NA_2 0 6.6452709208363170e-001
*
* Real pole n. 11
CS_11 NS_11 0 9.9999999999999998e-013
RS_11 NS_11 0 3.6187013423789601e+001
GS_11_2 0 NS_11 NA_2 0 6.6452709208363170e-001
*
* Real pole n. 12
CS_12 NS_12 0 9.9999999999999998e-013
RS_12 NS_12 0 4.6620502512561899e+002
GS_12_2 0 NS_12 NA_2 0 6.6452709208363170e-001
*
* Real pole n. 13
CS_13 NS_13 0 9.9999999999999998e-013
RS_13 NS_13 0 3.0454843143654548e+003
GS_13_2 0 NS_13 NA_2 0 6.6452709208363170e-001
*
* Real pole n. 14
CS_14 NS_14 0 9.9999999999999998e-013
RS_14 NS_14 0 4.2483511278785496e+004
GS_14_2 0 NS_14 NA_2 0 6.6452709208363170e-001
*
* Real pole n. 15
CS_15 NS_15 0 9.9999999999999998e-013
RS_15 NS_15 0 1.7479012563424539e+007
GS_15_2 0 NS_15 NA_2 0 6.6452709208363170e-001
*
* Real pole n. 16
CS_16 NS_16 0 9.9999999999999998e-013
RS_16 NS_16 0 7.6442948626474559e+007
GS_16_2 0 NS_16 NA_2 0 6.6452709208363170e-001
*
* Real pole n. 17
CS_17 NS_17 0 9.9999999999999998e-013
RS_17 NS_17 0 2.9502412466187273e+000
GS_17_3 0 NS_17 NA_3 0 6.6452709208363170e-001
*
* Real pole n. 18
CS_18 NS_18 0 9.9999999999999998e-013
RS_18 NS_18 0 9.7963963778649585e+000
GS_18_3 0 NS_18 NA_3 0 6.6452709208363170e-001
*
* Real pole n. 19
CS_19 NS_19 0 9.9999999999999998e-013
RS_19 NS_19 0 3.6187013423789601e+001
GS_19_3 0 NS_19 NA_3 0 6.6452709208363170e-001
*
* Real pole n. 20
CS_20 NS_20 0 9.9999999999999998e-013
RS_20 NS_20 0 4.6620502512561899e+002
GS_20_3 0 NS_20 NA_3 0 6.6452709208363170e-001
*
* Real pole n. 21
CS_21 NS_21 0 9.9999999999999998e-013
RS_21 NS_21 0 3.0454843143654548e+003
GS_21_3 0 NS_21 NA_3 0 6.6452709208363170e-001
*
* Real pole n. 22
CS_22 NS_22 0 9.9999999999999998e-013
RS_22 NS_22 0 4.2483511278785496e+004
GS_22_3 0 NS_22 NA_3 0 6.6452709208363170e-001
*
* Real pole n. 23
CS_23 NS_23 0 9.9999999999999998e-013
RS_23 NS_23 0 1.7479012563424539e+007
GS_23_3 0 NS_23 NA_3 0 6.6452709208363170e-001
*
* Real pole n. 24
CS_24 NS_24 0 9.9999999999999998e-013
RS_24 NS_24 0 7.6442948626474559e+007
GS_24_3 0 NS_24 NA_3 0 6.6452709208363170e-001
*
******************************


.ends
*******************
* End of subcircuit
*******************
.ends z90b_ondie_decoupling_perdq

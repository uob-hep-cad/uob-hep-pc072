* On-die Decoupling circuit for Z90B (VDDQ to VSSQ)
* Includes VDDQ-VSSQ decoupling for all signals (full die) including DQ0-15, LDQS_t/c, UDQS_t/c, UDM or LDM.
* This subcircuit should be added across the IBIS DQ, DM or DQS models' [Pullup Reference] and [Pulldown Reference]
* nodes as in the following Spice example:

******************************************************************************************************
*x_decouple vddq_die vcc_die vssq_die gnd z90b_ondie_decoupling_alldq

*b_dq1 vccq_die vssq_die PAD_DQ1 IN_DQ1 ENOUT RCVR_OUT_DQ1 vccq_die vssq_die
*+ file='z90b.ibs' model='DQ_34_2666' typ=typ power=off buffer=3 interpol=1 ramp_fwf=2 ramp_rwf=2
*+ rm_tail_rwf=default rm_tail_fwf=default
*+ rm_dly_rwf=default rm_dly_fwf=default
******************************************************************************************************


.subckt z90b_ondie_decoupling_alldq vddq_die vcc_die vssq_die ref
x1 vddq_die ref vcc_die ref vssq_die ref z90b_cfat_alldq


**********************************************************
** STATE-SPACE REALIZATION               
** IN SPICE LANGUAGE
** This file is automatically generated  
**********************************************************
** Created: 05-Apr-2018 by IdEM R2012 (8.0.6)
**********************************************************


**********************************************************
* NOTE:
* a_i  --> input node associated to the port i 
* b_i  --> reference node associated to the port i 
**********************************************************

***********************************
* Interface (ports specification) *
***********************************
.subckt z90b_cfat_alldq
+  a_1 b_1 
+  a_2 b_2 
+  a_3 b_3 
***********************************


******************************************
* Main circuit connected to output nodes *
******************************************

* Port 1
VI_1 a_1 NI_1 0
RI_1 NI_1 b_1 5.0000000000000000e+001
GC_1_1 b_1 NI_1 NS_1 0 1.7708196700277176e-003
GC_1_2 b_1 NI_1 NS_2 0 1.2892640209931625e-003
GC_1_3 b_1 NI_1 NS_3 0 1.0154872774493493e-003
GC_1_4 b_1 NI_1 NS_4 0 1.7324201084798801e-002
GC_1_5 b_1 NI_1 NS_5 0 5.2697455471491734e-005
GC_1_6 b_1 NI_1 NS_6 0 2.4830974709410387e-008
GC_1_7 b_1 NI_1 NS_7 0 1.3774272128278802e-006
GC_1_8 b_1 NI_1 NS_8 0 -1.6838460862776780e-013
GC_1_9 b_1 NI_1 NS_9 0 1.8210694709212458e-003
GC_1_10 b_1 NI_1 NS_10 0 1.2587484794872768e-003
GC_1_11 b_1 NI_1 NS_11 0 1.1182665786244213e-003
GC_1_12 b_1 NI_1 NS_12 0 1.7340069944902982e-002
GC_1_13 b_1 NI_1 NS_13 0 -1.0369064999302146e-004
GC_1_14 b_1 NI_1 NS_14 0 -3.5729019163142852e-008
GC_1_15 b_1 NI_1 NS_15 0 7.8545033063023424e-009
GC_1_16 b_1 NI_1 NS_16 0 4.3046844923824344e-013
GC_1_17 b_1 NI_1 NS_17 0 1.7215056561649756e-003
GC_1_18 b_1 NI_1 NS_18 0 1.3161919038290686e-003
GC_1_19 b_1 NI_1 NS_19 0 1.0245284322989248e-003
GC_1_20 b_1 NI_1 NS_20 0 1.7306358957883756e-002
GC_1_21 b_1 NI_1 NS_21 0 5.1803140885846370e-005
GC_1_22 b_1 NI_1 NS_22 0 1.0538549757757638e-008
GC_1_23 b_1 NI_1 NS_23 0 -1.3849859391838608e-006
GC_1_24 b_1 NI_1 NS_24 0 -2.6208533534192509e-013
GD_1_1 b_1 NI_1 NA_1 0 -2.7880389819231011e-001
GD_1_2 b_1 NI_1 NA_2 0 3.9001553882602618e-003
GD_1_3 b_1 NI_1 NA_3 0 3.9187482718857471e-003
*
* Port 2
VI_2 a_2 NI_2 0
RI_2 NI_2 b_2 5.0000000000000000e+001
GC_2_1 b_2 NI_2 NS_1 0 1.8210694709212452e-003
GC_2_2 b_2 NI_2 NS_2 0 1.2587484794872774e-003
GC_2_3 b_2 NI_2 NS_3 0 1.1182665786244211e-003
GC_2_4 b_2 NI_2 NS_4 0 1.7340069944902982e-002
GC_2_5 b_2 NI_2 NS_5 0 -1.0369064999302146e-004
GC_2_6 b_2 NI_2 NS_6 0 -3.5729019163143632e-008
GC_2_7 b_2 NI_2 NS_7 0 7.8545033063023903e-009
GC_2_8 b_2 NI_2 NS_8 0 4.3046844923808623e-013
GC_2_9 b_2 NI_2 NS_9 0 2.3310723434625934e-003
GC_2_10 b_2 NI_2 NS_10 0 1.3206040686207137e-003
GC_2_11 b_2 NI_2 NS_11 0 1.2082850712507624e-003
GC_2_12 b_2 NI_2 NS_12 0 1.7397485219076598e-002
GC_2_13 b_2 NI_2 NS_13 0 2.0402975959599176e-004
GC_2_14 b_2 NI_2 NS_14 0 4.5023381889150381e-008
GC_2_15 b_2 NI_2 NS_15 0 1.4586809863432922e-008
GC_2_16 b_2 NI_2 NS_16 0 -1.1005953563204874e-012
GC_2_17 b_2 NI_2 NS_17 0 1.8724309315601994e-003
GC_2_18 b_2 NI_2 NS_18 0 1.2735025892468838e-003
GC_2_19 b_2 NI_2 NS_19 0 1.1166396470161306e-003
GC_2_20 b_2 NI_2 NS_20 0 1.7329208767845612e-002
GC_2_21 b_2 NI_2 NS_21 0 -1.0192949552772539e-004
GC_2_22 b_2 NI_2 NS_22 0 -9.5431710035375882e-009
GC_2_23 b_2 NI_2 NS_23 0 -2.2438416263119445e-008
GC_2_24 b_2 NI_2 NS_24 0 6.7012753499802763e-013
GD_2_1 b_2 NI_2 NA_1 0 3.9001553882602618e-003
GD_2_2 b_2 NI_2 NA_2 0 -2.7879322778352789e-001
GD_2_3 b_2 NI_2 NA_3 0 4.0151906251375156e-003
*
* Port 3
VI_3 a_3 NI_3 0
RI_3 NI_3 b_3 5.0000000000000000e+001
GC_3_1 b_3 NI_3 NS_1 0 1.7215056561649756e-003
GC_3_2 b_3 NI_3 NS_2 0 1.3161919038290689e-003
GC_3_3 b_3 NI_3 NS_3 0 1.0245284322989245e-003
GC_3_4 b_3 NI_3 NS_4 0 1.7306358957883756e-002
GC_3_5 b_3 NI_3 NS_5 0 5.1803140885846390e-005
GC_3_6 b_3 NI_3 NS_6 0 1.0538549757756266e-008
GC_3_7 b_3 NI_3 NS_7 0 -1.3849859391838608e-006
GC_3_8 b_3 NI_3 NS_8 0 -2.6208533534218646e-013
GC_3_9 b_3 NI_3 NS_9 0 1.8724309315601994e-003
GC_3_10 b_3 NI_3 NS_10 0 1.2735025892468834e-003
GC_3_11 b_3 NI_3 NS_11 0 1.1166396470161306e-003
GC_3_12 b_3 NI_3 NS_12 0 1.7329208767845612e-002
GC_3_13 b_3 NI_3 NS_13 0 -1.0192949552772539e-004
GC_3_14 b_3 NI_3 NS_14 0 -9.5431710035381738e-009
GC_3_15 b_3 NI_3 NS_15 0 -2.2438416263119409e-008
GC_3_16 b_3 NI_3 NS_16 0 6.7012753499792838e-013
GC_3_17 b_3 NI_3 NS_17 0 1.8148358983513329e-003
GC_3_18 b_3 NI_3 NS_18 0 1.2955264578827608e-003
GC_3_19 b_3 NI_3 NS_19 0 1.0432266891081717e-003
GC_3_20 b_3 NI_3 NS_20 0 1.7286664617960350e-002
GC_3_21 b_3 NI_3 NS_21 0 5.0922247812203637e-005
GC_3_22 b_3 NI_3 NS_22 0 -1.3487518021214958e-009
GC_3_23 b_3 NI_3 NS_23 0 1.4071502256171362e-006
GC_3_24 b_3 NI_3 NS_24 0 -4.0804303737817002e-013
GD_3_1 b_3 NI_3 NA_1 0 3.9187482718857471e-003
GD_3_2 b_3 NI_3 NA_2 0 4.0151906251375156e-003
GD_3_3 b_3 NI_3 NA_3 0 -2.7882377530156416e-001
*
******************************************


********************************
* Synthesis of impinging waves *
********************************

* Impinging wave, port 1
RA_1 NA_1 0 3.5355339059327378e+000
FA_1 0 NA_1 VI_1 1.0
GA_1 0 NA_1 a_1 b_1 2.0000000000000000e-002
*
* Impinging wave, port 2
RA_2 NA_2 0 3.5355339059327378e+000
FA_2 0 NA_2 VI_2 1.0
GA_2 0 NA_2 a_2 b_2 2.0000000000000000e-002
*
* Impinging wave, port 3
RA_3 NA_3 0 3.5355339059327378e+000
FA_3 0 NA_3 VI_3 1.0
GA_3 0 NA_3 a_3 b_3 2.0000000000000000e-002
*
********************************


***************************************
* Synthesis of real and complex poles *
***************************************

* Real pole n. 1
CS_1 NS_1 0 9.9999999999999998e-013
RS_1 NS_1 0 9.7743856390692017e+000
GS_1_1 0 NS_1 NA_1 0 1.8408380925316373e-001
*
* Real pole n. 2
CS_2 NS_2 0 9.9999999999999998e-013
RS_2 NS_2 0 1.8515660105636602e+001
GS_2_1 0 NS_2 NA_1 0 1.8408380925316373e-001
*
* Real pole n. 3
CS_3 NS_3 0 9.9999999999999998e-013
RS_3 NS_3 0 3.8375109793817167e+001
GS_3_1 0 NS_3 NA_1 0 1.8408380925316373e-001
*
* Real pole n. 4
CS_4 NS_4 0 9.9999999999999998e-013
RS_4 NS_4 0 5.3029173403440033e+001
GS_4_1 0 NS_4 NA_1 0 1.8408380925316373e-001
*
* Real pole n. 5
CS_5 NS_5 0 9.9999999999999998e-013
RS_5 NS_5 0 9.7012921799809919e+003
GS_5_1 0 NS_5 NA_1 0 1.8408380925316373e-001
*
* Real pole n. 6
CS_6 NS_6 0 9.9999999999999998e-013
RS_6 NS_6 0 2.3964311160719226e+004
GS_6_1 0 NS_6 NA_1 0 1.8408380925316373e-001
*
* Real pole n. 7
CS_7 NS_7 0 9.9999999999999998e-013
RS_7 NS_7 0 2.4159751582315346e+005
GS_7_1 0 NS_7 NA_1 0 1.8408380925316373e-001
*
* Real pole n. 8
CS_8 NS_8 0 9.9999999999999998e-013
RS_8 NS_8 0 2.0999748010100037e+010
GS_8_1 0 NS_8 NA_1 0 1.8408380925316373e-001
*
* Real pole n. 9
CS_9 NS_9 0 9.9999999999999998e-013
RS_9 NS_9 0 9.7743856390692017e+000
GS_9_2 0 NS_9 NA_2 0 1.8408380925316373e-001
*
* Real pole n. 10
CS_10 NS_10 0 9.9999999999999998e-013
RS_10 NS_10 0 1.8515660105636602e+001
GS_10_2 0 NS_10 NA_2 0 1.8408380925316373e-001
*
* Real pole n. 11
CS_11 NS_11 0 9.9999999999999998e-013
RS_11 NS_11 0 3.8375109793817167e+001
GS_11_2 0 NS_11 NA_2 0 1.8408380925316373e-001
*
* Real pole n. 12
CS_12 NS_12 0 9.9999999999999998e-013
RS_12 NS_12 0 5.3029173403440033e+001
GS_12_2 0 NS_12 NA_2 0 1.8408380925316373e-001
*
* Real pole n. 13
CS_13 NS_13 0 9.9999999999999998e-013
RS_13 NS_13 0 9.7012921799809919e+003
GS_13_2 0 NS_13 NA_2 0 1.8408380925316373e-001
*
* Real pole n. 14
CS_14 NS_14 0 9.9999999999999998e-013
RS_14 NS_14 0 2.3964311160719226e+004
GS_14_2 0 NS_14 NA_2 0 1.8408380925316373e-001
*
* Real pole n. 15
CS_15 NS_15 0 9.9999999999999998e-013
RS_15 NS_15 0 2.4159751582315346e+005
GS_15_2 0 NS_15 NA_2 0 1.8408380925316373e-001
*
* Real pole n. 16
CS_16 NS_16 0 9.9999999999999998e-013
RS_16 NS_16 0 2.0999748010100037e+010
GS_16_2 0 NS_16 NA_2 0 1.8408380925316373e-001
*
* Real pole n. 17
CS_17 NS_17 0 9.9999999999999998e-013
RS_17 NS_17 0 9.7743856390692017e+000
GS_17_3 0 NS_17 NA_3 0 1.8408380925316373e-001
*
* Real pole n. 18
CS_18 NS_18 0 9.9999999999999998e-013
RS_18 NS_18 0 1.8515660105636602e+001
GS_18_3 0 NS_18 NA_3 0 1.8408380925316373e-001
*
* Real pole n. 19
CS_19 NS_19 0 9.9999999999999998e-013
RS_19 NS_19 0 3.8375109793817167e+001
GS_19_3 0 NS_19 NA_3 0 1.8408380925316373e-001
*
* Real pole n. 20
CS_20 NS_20 0 9.9999999999999998e-013
RS_20 NS_20 0 5.3029173403440033e+001
GS_20_3 0 NS_20 NA_3 0 1.8408380925316373e-001
*
* Real pole n. 21
CS_21 NS_21 0 9.9999999999999998e-013
RS_21 NS_21 0 9.7012921799809919e+003
GS_21_3 0 NS_21 NA_3 0 1.8408380925316373e-001
*
* Real pole n. 22
CS_22 NS_22 0 9.9999999999999998e-013
RS_22 NS_22 0 2.3964311160719226e+004
GS_22_3 0 NS_22 NA_3 0 1.8408380925316373e-001
*
* Real pole n. 23
CS_23 NS_23 0 9.9999999999999998e-013
RS_23 NS_23 0 2.4159751582315346e+005
GS_23_3 0 NS_23 NA_3 0 1.8408380925316373e-001
*
* Real pole n. 24
CS_24 NS_24 0 9.9999999999999998e-013
RS_24 NS_24 0 2.0999748010100037e+010
GS_24_3 0 NS_24 NA_3 0 1.8408380925316373e-001
*
******************************


.ends  z90b_cfat_alldq
*******************
* End of subcircuit
*******************
.ends  z90b_ondie_decoupling_alldq
